module ALU_tb();

    reg [31:0] Rtypr;
    reg [31:0] Itype;
    wire [31:0] Y;
    reg [31:0] Rtype,Itype;
    
    ALU F1(Rtype,Itype,Y);
    
    initial 
        begin
        Rtype = 32'b00000000000000000000000000000000;
        Itype = 32'b00000000000000000000000000000000;
        #10 Rtype = 32'b00000000000000000000000000000000;
        #10 Rtype = 32'b00000100000000000000000000000000;
        #10 Rtype = 32'b00001000000000000000000000000000;
        #10 Rtype = 32'b00001100000000000000000000000000;
        #10 Rtype = 32'b00010000000000000000000000000000;
        #10 Rtype = 32'b00010100000000000000000000000000;
        #10 Rtype = 32'b00011000000000000000000000000000;
        #10 Rtype = 32'b00101000000000000000000000000000;
        #10 Rtype = 32'b00101100000000000000000000000000; 
        #10 $stop;        
        end
    
endmodule
